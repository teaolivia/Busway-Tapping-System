-- controller