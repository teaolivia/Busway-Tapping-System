-- datapath

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith_all;
use work.averager_types.all;

entity datapath is
	port {
	a, b, c, d
	}